

library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use work.vga_package.all;

package Skyscrapers_Puzzle_Sprites is

	-- Game sprites:	
	type sprite_digits is array( 0 to 2024) of color_type; -- (24 * 24) color_type
	
CONSTANT zero_sprite: sprite_digits := (
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"555",X"777",X"777",X"777",X"777",X"777",X"555",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"BBB",X"BBB",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"DDD",X"DDD",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"FFF",X"FFF",X"FFF",X"DDD",X"777",X"333",X"333",X"111",X"333",X"333",X"555",X"999",X"FFF",X"FFF",X"FFF",X"DDD",X"111",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"FFF",X"777",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"BBB",X"FFF",X"DDD",X"DDD",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"FFF",X"777",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"BBB",X"FFF",X"DDD",X"DDD",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"FFF",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"FFF",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"DDD",X"DDD",X"FFF",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"777",X"FFF",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"FFF",X"999",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"555",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"555",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"555",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"555",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"111",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"FFF",X"777",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"BBB",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"FFF",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"FFF",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"FFF",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"FFF",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"777",X"FFF",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"FFF",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"777",X"FFF",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"DDD",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"FFF",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"FFF",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"FFF",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"FFF",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"FFF",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"FFF",X"999",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"DDD",X"FFF",X"111",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"FFF",X"777",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"555",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"333",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"555",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"333",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"FFF",X"BBB",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"FFF",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"999",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"FFF",X"FFF",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"DDD",X"DDD",X"FFF",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"DDD",X"FFF",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"FFF",X"FFF",X"999",X"999",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"DDD",X"FFF",X"BBB",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"FFF",X"FFF",X"999",X"999",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"DDD",X"FFF",X"BBB",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"DDD",X"FFF",X"FFF",X"FFF",X"999",X"777",X"777",X"555",X"555",X"555",X"777",X"BBB",X"FFF",X"FFF",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"777",X"DDD",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"BBB",X"BBB",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"333",X"333",X"555",X"555",X"555",X"333",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000"
);

CONSTANT one_sprite: sprite_digits := (
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"111",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"DDD",X"DDD",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"DDD",X"FFF",X"FFF",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"FFF",X"777",X"777",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"FFF",X"777",X"777",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"FFF",X"DDD",X"333",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"BBB",X"BBB",X"FFF",X"DDD",X"DDD",X"111",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"DDD",X"FFF",X"FFF",X"999",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"FFF",X"FFF",X"777",X"777",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"FFF",X"FFF",X"777",X"777",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"999",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"777",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000"
);

CONSTANT two_sprite: sprite_digits := (
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"555",X"777",X"777",X"777",X"777",X"777",X"777",X"555",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"999",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"999",X"999",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"BBB",X"FFF",X"FFF",X"FFF",X"DDD",X"999",X"999",X"555",X"333",X"111",X"111",X"333",X"555",X"555",X"777",X"DDD",X"FFF",X"FFF",X"FFF",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"BBB",X"FFF",X"FFF",X"FFF",X"DDD",X"999",X"999",X"555",X"333",X"111",X"111",X"333",X"555",X"555",X"777",X"DDD",X"FFF",X"FFF",X"FFF",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"999",X"999",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"999",X"FFF",X"FFF",X"333",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"BBB",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"FFF",X"FFF",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"FFF",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"FFF",X"FFF",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"DDD",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"555",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"DDD",X"DDD",X"FFF",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"DDD",X"111",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"DDD",X"111",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"FFF",X"FFF",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"FFF",X"FFF",X"FFF",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"FFF",X"FFF",X"333",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"FFF",X"FFF",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"FFF",X"FFF",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"FFF",X"333",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"FFF",X"FFF",X"FFF",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"FFF",X"DDD",X"DDD",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"999",X"FFF",X"DDD",X"111",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"999",X"FFF",X"DDD",X"111",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"BBB",X"FFF",X"FFF",X"BBB",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"FFF",X"FFF",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000"
);

CONSTANT three_sprite: sprite_digits := (
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"555",X"777",X"777",X"777",X"999",X"777",X"777",X"555",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"999",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"DDD",X"DDD",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"FFF",X"FFF",X"BBB",X"777",X"777",X"555",X"333",X"111",X"111",X"111",X"333",X"333",X"555",X"999",X"FFF",X"FFF",X"FFF",X"DDD",X"111",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"999",X"999",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"BBB",X"FFF",X"BBB",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"999",X"999",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"BBB",X"FFF",X"BBB",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"DDD",X"FFF",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"FFF",X"FFF",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"FFF",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"FFF",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"FFF",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"FFF",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"FFF",X"DDD",X"333",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"777",X"DDD",X"FFF",X"FFF",X"BBB",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"BBB",X"BBB",X"BBB",X"BBB",X"DDD",X"DDD",X"FFF",X"FFF",X"FFF",X"FFF",X"999",X"333",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"BBB",X"BBB",X"BBB",X"BBB",X"DDD",X"DDD",X"FFF",X"FFF",X"FFF",X"FFF",X"999",X"333",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"DDD",X"999",X"333",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"111",X"111",X"111",X"111",X"333",X"777",X"777",X"999",X"FFF",X"FFF",X"FFF",X"DDD",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"DDD",X"FFF",X"777",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"DDD",X"FFF",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"DDD",X"FFF",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"FFF",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"DDD",X"DDD",X"FFF",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"999",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"999",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"777",X"FFF",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"999",X"FFF",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"FFF",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"FFF",X"FFF",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"FFF",X"FFF",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"DDD",X"777",X"777",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"777",X"777",X"FFF",X"FFF",X"777",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"DDD",X"777",X"777",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"777",X"777",X"FFF",X"FFF",X"777",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"DDD",X"FFF",X"FFF",X"FFF",X"BBB",X"999",X"999",X"555",X"555",X"555",X"555",X"555",X"777",X"777",X"BBB",X"FFF",X"FFF",X"FFF",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"555",X"999",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"DDD",X"777",X"777",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"333",X"555",X"555",X"555",X"555",X"333",X"333",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000"
);

CONSTANT four_sprite: sprite_digits := (
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"DDD",X"FFF",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"FFF",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"FFF",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"FFF",X"999",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"333",X"FFF",X"DDD",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"DDD",X"DDD",X"FFF",X"333",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"FFF",X"FFF",X"777",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"FFF",X"BBB",X"BBB",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"FFF",X"BBB",X"BBB",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"FFF",X"DDD",X"111",X"111",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"FFF",X"FFF",X"999",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"DDD",X"DDD",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"DDD",X"FFF",X"111",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"111",X"DDD",X"FFF",X"111",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"999",X"999",X"FFF",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"FFF",X"FFF",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"FFF",X"DDD",X"DDD",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"333",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"FFF",X"333",X"333",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"777",X"777",X"FFF",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"333",X"FFF",X"FFF",X"BBB",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"111",X"DDD",X"FFF",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"FFF",X"FFF",X"FFF",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"FFF",X"FFF",X"FFF",X"FFF",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"DDD",X"777",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"FFF",X"FFF",X"FFF",X"DDD",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"555",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"FFF",X"FFF",X"FFF",X"DDD",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"BBB",X"555",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"BBB",X"BBB",X"FFF",X"111",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",
	X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000"
);

end package;